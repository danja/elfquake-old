.title KiCad schematic
U1 Net-_C2-Pad1_ Net-_R2-Pad1_ Net-_C1-Pad2_ Net-_C13-Pad1_ Net-_C3-Pad2_ Net-_C6-Pad1_ Net-_C6-Pad1_ Net-_RV1-Pad1_ Net-_RV1-Pad1_ Net-_C7-Pad2_ Net-_C14-Pad2_ Net-_C10-Pad2_ Net-_R12-Pad1_ Net-_D1-Pad1_ TL074
R3 Net-_C2-Pad1_ Net-_R2-Pad1_ 100k
R1 Net-_C1-Pad2_ 0 10M
R2 Net-_R2-Pad1_ 0 10k
SW1 +9V Net-_C13-Pad1_ NC_01 -9V Net-_C14-Pad2_ NC_02 SW_DPDT_x2
AE1 Net-_AE1-Pad1_ Antenna
C1 Net-_AE1-Pad1_ Net-_C1-Pad2_ 10n
C5 Net-_C4-Pad1_ 0 100n
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 100n
C3 Net-_C2-Pad2_ Net-_C3-Pad2_ 100n
R6 Net-_C2-Pad2_ 0 15k
R4 Net-_C2-Pad1_ Net-_C4-Pad1_ 33k
R5 Net-_C4-Pad1_ Net-_C3-Pad2_ 33k
C4 Net-_C4-Pad1_ 0 100n
C9 Net-_C8-Pad1_ 0 47n
C6 Net-_C6-Pad1_ Net-_C6-Pad2_ 47n
C7 Net-_C6-Pad2_ Net-_C7-Pad2_ 47n
R9 Net-_C6-Pad2_ 0 22k
R7 Net-_C6-Pad1_ Net-_C8-Pad1_ 22k
R8 Net-_C8-Pad1_ Net-_C7-Pad2_ 22k
C8 Net-_C8-Pad1_ 0 47n
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ 1N4148
D2 Net-_D2-Pad1_ Net-_D1-Pad1_ 1N4148
Q1 Net-_C12-Pad1_ Net-_D1-Pad2_ Net-_C13-Pad1_ 2N3904
Q2 Net-_C14-Pad2_ Net-_D2-Pad1_ Net-_C12-Pad1_ 2N3906
R15 Net-_C13-Pad1_ Net-_D1-Pad2_ 8k2
R16 Net-_D2-Pad1_ Net-_C14-Pad2_ 8k2
R12 Net-_R12-Pad1_ Net-_C12-Pad1_ 100k
R13 Net-_R12-Pad1_ Net-_C11-Pad1_ 1k5
R14 Net-_C11-Pad1_ 0 10k
C11 Net-_C11-Pad1_ 0 1u
C13 Net-_C13-Pad1_ 0 100u
C14 0 Net-_C14-Pad2_ 100u
C12 Net-_C12-Pad1_ Net-_C12-Pad2_ 100u
LS1 Net-_C12-Pad2_ 0 8
C10 Net-_C10-Pad1_ Net-_C10-Pad2_ 10u
R11 Net-_C10-Pad2_ 0 1M
RV1 Net-_RV1-Pad1_ Net-_C10-Pad1_ 0 100k
R10 Net-_C6-Pad2_ 0 22k
J1 Net-_AE1-Pad1_ Conn_01x01_Female
.end
